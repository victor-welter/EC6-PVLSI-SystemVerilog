module exe_02
(
    input logic btn_n_i,
	
    output logic led_n_o
);

assign led_n_o = btn_n_i;

endmodule